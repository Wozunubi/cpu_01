module datapath #(
  
) (
  input logic clk,
  
);



endmodule